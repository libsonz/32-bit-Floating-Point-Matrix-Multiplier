`timescale 1ns / 1ps

module multiplier_32bit_tb();

    // DUT signals
    reg [31:0] i_a, i_b;
    reg        i_vld;
    wire [31:0] o_res;
    wire        o_res_vld;
    wire        overflow;

    // Counters
    integer pass_count = 0;
    integer fail_count = 0;
    integer test_num = 0;

    // Instantiate DUT
    multiplier_32bit uut (
        .i_a(i_a),
        .i_b(i_b),
        .i_vld(i_vld),
        .o_res(o_res),
        .o_res_vld(o_res_vld),
        .overflow(overflow)
    );

    // Task to run a single test case
    task automatic run_test;
        input [31:0] a_val;
        input [31:0] b_val;
        input [31:0] expected;
        begin
            test_num = test_num + 1;
            i_a = a_val;
            i_b = b_val;
            i_vld = 1'b1;
            #1;
            i_vld = 1'b0;

            // Wait for output valid
            wait(o_res_vld === 1'b1);
            #1;
            
            $display("Test %0d:", test_num);
            $display("  Input A:   0x%08h", a_val);
            $display("  Input B:   0x%08h", b_val);
            $display("  Expected:  0x%08h", expected);
            $display("  Actual:    0x%08h", o_res);
            $display("  Overflow:  %b", overflow);

            if (o_res === expected) begin
                $display("  Result: PASS\n");
                pass_count = pass_count + 1;
            end else begin
                $display("  Result: FAIL\n");
                fail_count = fail_count + 1;
            end

            // Wait for o_res_vld to deassert before next test
            wait(o_res_vld === 1'b0);
            #1;
        end
    endtask

    // Hex values from scripts/floating_point.py output
    // Example:
    // // 2.0 * 3.0 = 6.0
    // run_test(32'h40000000, 32'h40400000, 32'h40c00000);

    initial begin
        $display("\nStarting multiplier_32bit testbench\n");

        // Test Cases generated by scripts/floating_point.py
        run_test(32'h40000000, 32'h40400000, 32'h40c00000); // 2.0 * 3.0 = 6.0
        run_test(32'hc0000000, 32'h40400000, 32'hc0c00000); // -2.0 * 3.0 = -6.0
        run_test(32'h00000000, 32'h42f6e979, 32'h00000000); // 0.0 * 123.456 = 0.0
        run_test(32'h7f800000, 32'h40000000, 32'h7f800000); // inf * 2.0 = inf
        run_test(32'h7f800000, 32'hc0000000, 32'hff800000); // inf * -2.0 = -inf
        run_test(32'h7fc00000, 32'h40000000, 32'h7fc00000); // nan * 2.0 = nan
        run_test(32'h7f800000, 32'h00000000, 32'h7fc00000); // inf * 0.0 = nan
        run_test(32'h3fc00000, 32'hc0880000, 32'hc0a70000); // 1.5 * -4.25 = -6.375
        run_test(32'h4123ae14, 32'hc0880000, 32'hc214b972); // 10.24 * -4.25 = -43.52
        run_test(32'h2f5c28f6, 32'hc1205e6e, 32'hbfe4c4f5); // 1e-9 * -10.88888888 = -1.08888889e-08

        $display("\nTestbench Complete");
        $display("Tests Run: %0d", test_num);
        $display("Passed:    %0d", pass_count);
        $display("Failed:    %0d", fail_count);

        if (fail_count == 0) $display("SUCCESS: All tests passed!");
        else                 $display("FAILURE: Some tests failed.");

        #10 $finish;
    end

    // Optional: VCD dump for waveform viewing
    initial begin
        $dumpfile("multiplier_32bit_tb.vcd");
        $dumpvars(0, multiplier_32bit_tb);
    end

endmodule
